`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/08/27 09:38:11
// Design Name: 
// Module Name: delimiter_check
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module delimiter_check(
            input           rst,                    //��λ�ź�
            input           clk_3M,                 //3Mʱ���ź�
            input           clk_6M,                 //6Mʱ���ź�
            input           data_in,                //��������
            input           frame_end,              //֡ĩβ�ź�
            output reg      M_frame,               //��֡��ʼ�ź�
            output reg      S_frame,               //��֡��ʼ�ź�
            output reg      E_frame,               //֡��ֹ�ź�
            output reg      E_delimit,             //�ֽ�������ź�
            output reg      E_length               //���ȴ����ź�
    );
    reg[4:0]        delimiter_counter=5'h0;
    reg[15:0]       delimiter_in=16'h0;
    wire            data;
	parameter      M_delimiter=16'b1100011100010101;  
    parameter      S_delimiter=16'b1010100011100011;  
    parameter      E_delimiter=4'b0011;
    
    
    assign data=data_in^clk_3M;
    
    always @(negedge clk_6M or negedge rst)begin
        if(rst==1'b0)begin
            delimiter_in<=16'h0;
            delimiter_counter<=5'h0;
        end else begin
            delimiter_in[0]<=data_in;
            delimiter_in[15:1]<=delimiter_in[14:0];
            delimiter_counter<=delimiter_counter+1;
        end
    end
    
    always @(*) begin
        if(rst==1'b0)begin
            M_frame<=1'b0;
            S_frame<=1'b0;
            E_frame<=1'b0;
            E_delimit<=1'b0;
            E_length<=1'b0;
        end else if(delimiter_counter==5'h4&&frame_end==1'b1)begin
            if(delimiter_in[3:0]==E_delimiter)begin
                M_frame<=1'b0;
                S_frame<=1'b0;
                E_frame<=1'b1;
                E_delimit<=1'b0;
                E_length<=1'b0;                
            end  else begin
                M_frame<=1'b0;
                S_frame<=1'b0;
                E_frame<=1'b0;
                E_delimit<=1'b0;            
                E_length<=1'b1;
            end
        end  else if(delimiter_counter==5'h11)begin
                if(delimiter_in==M_delimiter)begin
                    M_frame<=1'b1;
                    S_frame<=1'b0;
                    E_frame<=1'b0;
                    E_delimit<=1'b0;
                    E_length<=1'b0;
                end else if(delimiter_in==S_delimiter)begin
                    S_frame<=1'b1;
                    M_frame<=1'b0;
                    E_frame<=1'b0;
                    E_delimit<=1'b0;
                    E_length<=1'b0;                
                end else begin
                    S_frame<=1'b0;
                    M_frame<=1'b0;
                    E_frame<=1'b0;
                    E_delimit<=1'b1;
                    E_length<=1'b0;
                end
        end else begin
            M_frame<=M_frame;
            S_frame<=S_frame;
            E_frame<=E_frame;
            E_delimit<=1'b0;
            E_length<=E_length;            
        end
     end
     

    
    
    
endmodule
